module signExtend(i_data, o_data);
input   [15:0]  i_data;
output  [31:0]  o_data;

endmodule