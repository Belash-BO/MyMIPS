`timescale 1ns / 1ps

module Shifter_tb;

	parameter period = 128;

	reg [4:0]	SA;
	reg [1:0]	SRO;
	reg [31:0]	Data;
	wire[31:0]	Result;
	integer i;
	integer j;

	Shifter Shifter_tb (.SA(SA), .SRO(SRO), .Data(Data), .Result(Result));

	initial begin
		forever #(period/128) begin
			for (i = 0; i <= 3; i = i + 1) #32 SRO = i;
		end
	end
	
	initial begin
		SA = 31;
		forever #(period/4) begin
			for (j = 0; j <= 31; j = j + 1) #1 SA = j;
		end
	end

	initial begin
		forever #(period/512) Data = $random;
	end

	initial #5000 $stop;
endmodule
